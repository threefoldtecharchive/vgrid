module model

// TODO: farm struct
