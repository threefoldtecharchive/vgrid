module model

// TODO: contract struct
